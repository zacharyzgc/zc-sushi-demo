/*
 * Copyright (c) 2024 ZC
 * SPDX-License-Identifier: Apache-2.0
 */


module tt_um_sushi_demo (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);
//  |-----------H_DISPLAY-----------|-----H_FRONT-----|-----H_SYNC-----|-----H_BACK-----|

  // horizontal constants
  parameter H_DISPLAY       = 640; // horizontal display width
  parameter H_BACK          =  48; // horizontal left border (back porch)
  parameter H_FRONT         =  16; // horizontal right border (front porch)
  parameter H_SYNC          =  96; // horizontal sync width
  // vertical constants
  parameter V_DISPLAY       = 480; // vertical display height
  parameter V_TOP           =  33; // vertical top border
  parameter V_BOTTOM        =  10; // vertical bottom border
  parameter V_SYNC          =   2; // vertical sync # lines
  // derived constants
  parameter H_SYNC_START    = H_DISPLAY + H_FRONT;
  parameter H_SYNC_END      = H_DISPLAY + H_FRONT + H_SYNC - 1;
  parameter H_MAX           = H_DISPLAY + H_BACK + H_FRONT + H_SYNC - 1;
  parameter V_SYNC_START    = V_DISPLAY + V_BOTTOM;
  parameter V_SYNC_END      = V_DISPLAY + V_BOTTOM + V_SYNC - 1;
  parameter V_MAX           = V_DISPLAY + V_TOP + V_BOTTOM + V_SYNC - 1;
  //sprite position
  parameter SPRITE_X_START = 100;
  parameter SPRITE_Y_START = 100;
  parameter SPRITE_WIDTH = 33*8;
  parameter SPRITE_HEIGHT = 19*8;

  //sprite frames
    
  reg [1:0] sushi_run_0 [18:0] [32:0]; //33x19 sprite [y][x]

  always @(*) begin
  sushi_run_0[0][0] = 2'b00;
  sushi_run_0[0][1] = 2'b00;
  sushi_run_0[0][2] = 2'b00;
  sushi_run_0[0][3] = 2'b00;
  sushi_run_0[0][4] = 2'b00;
  sushi_run_0[0][5] = 2'b00;
  sushi_run_0[0][6] = 2'b00;
  sushi_run_0[0][7] = 2'b00;
  sushi_run_0[0][8] = 2'b00;
  sushi_run_0[0][9] = 2'b00;
  sushi_run_0[0][10] = 2'b00;
  sushi_run_0[0][11] = 2'b00;
  sushi_run_0[0][12] = 2'b00;
  sushi_run_0[0][13] = 2'b00;
  sushi_run_0[0][14] = 2'b00;
  sushi_run_0[0][15] = 2'b00;
  sushi_run_0[0][16] = 2'b00;
  sushi_run_0[0][17] = 2'b00;
  sushi_run_0[0][18] = 2'b00;
  sushi_run_0[0][19] = 2'b00;
  sushi_run_0[0][20] = 2'b00;
  sushi_run_0[0][21] = 2'b00;
  sushi_run_0[0][22] = 2'b01;
  sushi_run_0[0][23] = 2'b01;
  sushi_run_0[0][24] = 2'b01;
  sushi_run_0[0][25] = 2'b01;
  sushi_run_0[0][26] = 2'b01;
  sushi_run_0[0][27] = 2'b01;
  sushi_run_0[0][28] = 2'b00;
  sushi_run_0[0][29] = 2'b00;
  sushi_run_0[0][30] = 2'b00;
  sushi_run_0[0][31] = 2'b00;
  sushi_run_0[0][32] = 2'b00;
  sushi_run_0[1][0] = 2'b00;
  sushi_run_0[1][1] = 2'b00;
  sushi_run_0[1][2] = 2'b00;
  sushi_run_0[1][3] = 2'b00;
  sushi_run_0[1][4] = 2'b00;
  sushi_run_0[1][5] = 2'b00;
  sushi_run_0[1][6] = 2'b00;
  sushi_run_0[1][7] = 2'b00;
  sushi_run_0[1][8] = 2'b00;
  sushi_run_0[1][9] = 2'b00;
  sushi_run_0[1][10] = 2'b00;
  sushi_run_0[1][11] = 2'b00;
  sushi_run_0[1][12] = 2'b00;
  sushi_run_0[1][13] = 2'b00;
  sushi_run_0[1][14] = 2'b00;
  sushi_run_0[1][15] = 2'b00;
  sushi_run_0[1][16] = 2'b00;
  sushi_run_0[1][17] = 2'b00;
  sushi_run_0[1][18] = 2'b00;
  sushi_run_0[1][19] = 2'b00;
  sushi_run_0[1][20] = 2'b00;
  sushi_run_0[1][21] = 2'b01;
  sushi_run_0[1][22] = 2'b01;
  sushi_run_0[1][23] = 2'b11;
  sushi_run_0[1][24] = 2'b10;
  sushi_run_0[1][25] = 2'b10;
  sushi_run_0[1][26] = 2'b10;
  sushi_run_0[1][27] = 2'b01;
  sushi_run_0[1][28] = 2'b01;
  sushi_run_0[1][29] = 2'b00;
  sushi_run_0[1][30] = 2'b00;
  sushi_run_0[1][31] = 2'b00;
  sushi_run_0[1][32] = 2'b00;
  sushi_run_0[2][0] = 2'b00;
  sushi_run_0[2][1] = 2'b00;
  sushi_run_0[2][2] = 2'b00;
  sushi_run_0[2][3] = 2'b00;
  sushi_run_0[2][4] = 2'b00;
  sushi_run_0[2][5] = 2'b00;
  sushi_run_0[2][6] = 2'b00;
  sushi_run_0[2][7] = 2'b00;
  sushi_run_0[2][8] = 2'b00;
  sushi_run_0[2][9] = 2'b00;
  sushi_run_0[2][10] = 2'b00;
  sushi_run_0[2][11] = 2'b00;
  sushi_run_0[2][12] = 2'b00;
  sushi_run_0[2][13] = 2'b00;
  sushi_run_0[2][14] = 2'b00;
  sushi_run_0[2][15] = 2'b00;
  sushi_run_0[2][16] = 2'b00;
  sushi_run_0[2][17] = 2'b00;
  sushi_run_0[2][18] = 2'b00;
  sushi_run_0[2][19] = 2'b00;
  sushi_run_0[2][20] = 2'b01;
  sushi_run_0[2][21] = 2'b01;
  sushi_run_0[2][22] = 2'b11;
  sushi_run_0[2][23] = 2'b10;
  sushi_run_0[2][24] = 2'b10;
  sushi_run_0[2][25] = 2'b10;
  sushi_run_0[2][26] = 2'b10;
  sushi_run_0[2][27] = 2'b10;
  sushi_run_0[2][28] = 2'b01;
  sushi_run_0[2][29] = 2'b01;
  sushi_run_0[2][30] = 2'b00;
  sushi_run_0[2][31] = 2'b00;
  sushi_run_0[2][32] = 2'b00;
  sushi_run_0[3][0] = 2'b00;
  sushi_run_0[3][1] = 2'b00;
  sushi_run_0[3][2] = 2'b00;
  sushi_run_0[3][3] = 2'b00;
  sushi_run_0[3][4] = 2'b00;
  sushi_run_0[3][5] = 2'b00;
  sushi_run_0[3][6] = 2'b00;
  sushi_run_0[3][7] = 2'b00;
  sushi_run_0[3][8] = 2'b00;
  sushi_run_0[3][9] = 2'b00;
  sushi_run_0[3][10] = 2'b00;
  sushi_run_0[3][11] = 2'b00;
  sushi_run_0[3][12] = 2'b00;
  sushi_run_0[3][13] = 2'b00;
  sushi_run_0[3][14] = 2'b00;
  sushi_run_0[3][15] = 2'b00;
  sushi_run_0[3][16] = 2'b00;
  sushi_run_0[3][17] = 2'b00;
  sushi_run_0[3][18] = 2'b00;
  sushi_run_0[3][19] = 2'b00;
  sushi_run_0[3][20] = 2'b01;
  sushi_run_0[3][21] = 2'b11;
  sushi_run_0[3][22] = 2'b10;
  sushi_run_0[3][23] = 2'b10;
  sushi_run_0[3][24] = 2'b10;
  sushi_run_0[3][25] = 2'b10;
  sushi_run_0[3][26] = 2'b10;
  sushi_run_0[3][27] = 2'b10;
  sushi_run_0[3][28] = 2'b10;
  sushi_run_0[3][29] = 2'b01;
  sushi_run_0[3][30] = 2'b00;
  sushi_run_0[3][31] = 2'b00;
  sushi_run_0[3][32] = 2'b00;
  sushi_run_0[4][0] = 2'b01;
  sushi_run_0[4][1] = 2'b01;
  sushi_run_0[4][2] = 2'b00;
  sushi_run_0[4][3] = 2'b00;
  sushi_run_0[4][4] = 2'b00;
  sushi_run_0[4][5] = 2'b00;
  sushi_run_0[4][6] = 2'b00;
  sushi_run_0[4][7] = 2'b00;
  sushi_run_0[4][8] = 2'b00;
  sushi_run_0[4][9] = 2'b00;
  sushi_run_0[4][10] = 2'b00;
  sushi_run_0[4][11] = 2'b00;
  sushi_run_0[4][12] = 2'b00;
  sushi_run_0[4][13] = 2'b00;
  sushi_run_0[4][14] = 2'b00;
  sushi_run_0[4][15] = 2'b00;
  sushi_run_0[4][16] = 2'b00;
  sushi_run_0[4][17] = 2'b00;
  sushi_run_0[4][18] = 2'b01;
  sushi_run_0[4][19] = 2'b01;
  sushi_run_0[4][20] = 2'b11;
  sushi_run_0[4][21] = 2'b10;
  sushi_run_0[4][22] = 2'b10;
  sushi_run_0[4][23] = 2'b10;
  sushi_run_0[4][24] = 2'b10;
  sushi_run_0[4][25] = 2'b10;
  sushi_run_0[4][26] = 2'b01;
  sushi_run_0[4][27] = 2'b01;
  sushi_run_0[4][28] = 2'b10;
  sushi_run_0[4][29] = 2'b01;
  sushi_run_0[4][30] = 2'b01;
  sushi_run_0[4][31] = 2'b00;
  sushi_run_0[4][32] = 2'b00;
  sushi_run_0[5][0] = 2'b01;
  sushi_run_0[5][1] = 2'b01;
  sushi_run_0[5][2] = 2'b01;
  sushi_run_0[5][3] = 2'b00;
  sushi_run_0[5][4] = 2'b00;
  sushi_run_0[5][5] = 2'b00;
  sushi_run_0[5][6] = 2'b00;
  sushi_run_0[5][7] = 2'b00;
  sushi_run_0[5][8] = 2'b00;
  sushi_run_0[5][9] = 2'b00;
  sushi_run_0[5][10] = 2'b00;
  sushi_run_0[5][11] = 2'b00;
  sushi_run_0[5][12] = 2'b00;
  sushi_run_0[5][13] = 2'b00;
  sushi_run_0[5][14] = 2'b00;
  sushi_run_0[5][15] = 2'b00;
  sushi_run_0[5][16] = 2'b00;
  sushi_run_0[5][17] = 2'b00;
  sushi_run_0[5][18] = 2'b01;
  sushi_run_0[5][19] = 2'b11;
  sushi_run_0[5][20] = 2'b11;
  sushi_run_0[5][21] = 2'b10;
  sushi_run_0[5][22] = 2'b10;
  sushi_run_0[5][23] = 2'b10;
  sushi_run_0[5][24] = 2'b10;
  sushi_run_0[5][25] = 2'b10;
  sushi_run_0[5][26] = 2'b10;
  sushi_run_0[5][27] = 2'b01;
  sushi_run_0[5][28] = 2'b01;
  sushi_run_0[5][29] = 2'b10;
  sushi_run_0[5][30] = 2'b01;
  sushi_run_0[5][31] = 2'b00;
  sushi_run_0[5][32] = 2'b00;
  sushi_run_0[6][0] = 2'b01;
  sushi_run_0[6][1] = 2'b01;
  sushi_run_0[6][2] = 2'b01;
  sushi_run_0[6][3] = 2'b01;
  sushi_run_0[6][4] = 2'b00;
  sushi_run_0[6][5] = 2'b00;
  sushi_run_0[6][6] = 2'b00;
  sushi_run_0[6][7] = 2'b00;
  sushi_run_0[6][8] = 2'b00;
  sushi_run_0[6][9] = 2'b00;
  sushi_run_0[6][10] = 2'b00;
  sushi_run_0[6][11] = 2'b00;
  sushi_run_0[6][12] = 2'b00;
  sushi_run_0[6][13] = 2'b00;
  sushi_run_0[6][14] = 2'b00;
  sushi_run_0[6][15] = 2'b00;
  sushi_run_0[6][16] = 2'b00;
  sushi_run_0[6][17] = 2'b00;
  sushi_run_0[6][18] = 2'b01;
  sushi_run_0[6][19] = 2'b11;
  sushi_run_0[6][20] = 2'b10;
  sushi_run_0[6][21] = 2'b10;
  sushi_run_0[6][22] = 2'b10;
  sushi_run_0[6][23] = 2'b10;
  sushi_run_0[6][24] = 2'b01;
  sushi_run_0[6][25] = 2'b10;
  sushi_run_0[6][26] = 2'b10;
  sushi_run_0[6][27] = 2'b01;
  sushi_run_0[6][28] = 2'b01;
  sushi_run_0[6][29] = 2'b10;
  sushi_run_0[6][30] = 2'b01;
  sushi_run_0[6][31] = 2'b01;
  sushi_run_0[6][32] = 2'b01;
  sushi_run_0[7][0] = 2'b00;
  sushi_run_0[7][1] = 2'b01;
  sushi_run_0[7][2] = 2'b10;
  sushi_run_0[7][3] = 2'b01;
  sushi_run_0[7][4] = 2'b00;
  sushi_run_0[7][5] = 2'b00;
  sushi_run_0[7][6] = 2'b00;
  sushi_run_0[7][7] = 2'b00;
  sushi_run_0[7][8] = 2'b00;
  sushi_run_0[7][9] = 2'b00;
  sushi_run_0[7][10] = 2'b00;
  sushi_run_0[7][11] = 2'b00;
  sushi_run_0[7][12] = 2'b00;
  sushi_run_0[7][13] = 2'b00;
  sushi_run_0[7][14] = 2'b00;
  sushi_run_0[7][15] = 2'b01;
  sushi_run_0[7][16] = 2'b01;
  sushi_run_0[7][17] = 2'b01;
  sushi_run_0[7][18] = 2'b01;
  sushi_run_0[7][19] = 2'b11;
  sushi_run_0[7][20] = 2'b10;
  sushi_run_0[7][21] = 2'b10;
  sushi_run_0[7][22] = 2'b10;
  sushi_run_0[7][23] = 2'b01;
  sushi_run_0[7][24] = 2'b01;
  sushi_run_0[7][25] = 2'b10;
  sushi_run_0[7][26] = 2'b10;
  sushi_run_0[7][27] = 2'b10;
  sushi_run_0[7][28] = 2'b10;
  sushi_run_0[7][29] = 2'b10;
  sushi_run_0[7][30] = 2'b10;
  sushi_run_0[7][31] = 2'b10;
  sushi_run_0[7][32] = 2'b01;
  sushi_run_0[8][0] = 2'b00;
  sushi_run_0[8][1] = 2'b01;
  sushi_run_0[8][2] = 2'b10;
  sushi_run_0[8][3] = 2'b01;
  sushi_run_0[8][4] = 2'b01;
  sushi_run_0[8][5] = 2'b01;
  sushi_run_0[8][6] = 2'b00;
  sushi_run_0[8][7] = 2'b01;
  sushi_run_0[8][8] = 2'b01;
  sushi_run_0[8][9] = 2'b01;
  sushi_run_0[8][10] = 2'b01;
  sushi_run_0[8][11] = 2'b01;
  sushi_run_0[8][12] = 2'b01;
  sushi_run_0[8][13] = 2'b01;
  sushi_run_0[8][14] = 2'b01;
  sushi_run_0[8][15] = 2'b01;
  sushi_run_0[8][16] = 2'b10;
  sushi_run_0[8][17] = 2'b11;
  sushi_run_0[8][18] = 2'b01;
  sushi_run_0[8][19] = 2'b01;
  sushi_run_0[8][20] = 2'b10;
  sushi_run_0[8][21] = 2'b10;
  sushi_run_0[8][22] = 2'b10;
  sushi_run_0[8][23] = 2'b01;
  sushi_run_0[8][24] = 2'b10;
  sushi_run_0[8][25] = 2'b10;
  sushi_run_0[8][26] = 2'b10;
  sushi_run_0[8][27] = 2'b10;
  sushi_run_0[8][28] = 2'b10;
  sushi_run_0[8][29] = 2'b10;
  sushi_run_0[8][30] = 2'b10;
  sushi_run_0[8][31] = 2'b01;
  sushi_run_0[8][32] = 2'b01;
  sushi_run_0[9][0] = 2'b00;
  sushi_run_0[9][1] = 2'b01;
  sushi_run_0[9][2] = 2'b01;
  sushi_run_0[9][3] = 2'b10;
  sushi_run_0[9][4] = 2'b10;
  sushi_run_0[9][5] = 2'b01;
  sushi_run_0[9][6] = 2'b01;
  sushi_run_0[9][7] = 2'b01;
  sushi_run_0[9][8] = 2'b10;
  sushi_run_0[9][9] = 2'b10;
  sushi_run_0[9][10] = 2'b10;
  sushi_run_0[9][11] = 2'b10;
  sushi_run_0[9][12] = 2'b10;
  sushi_run_0[9][13] = 2'b10;
  sushi_run_0[9][14] = 2'b10;
  sushi_run_0[9][15] = 2'b10;
  sushi_run_0[9][16] = 2'b10;
  sushi_run_0[9][17] = 2'b11;
  sushi_run_0[9][18] = 2'b10;
  sushi_run_0[9][19] = 2'b01;
  sushi_run_0[9][20] = 2'b01;
  sushi_run_0[9][21] = 2'b01;
  sushi_run_0[9][22] = 2'b01;
  sushi_run_0[9][23] = 2'b01;
  sushi_run_0[9][24] = 2'b10;
  sushi_run_0[9][25] = 2'b10;
  sushi_run_0[9][26] = 2'b10;
  sushi_run_0[9][27] = 2'b10;
  sushi_run_0[9][28] = 2'b10;
  sushi_run_0[9][29] = 2'b10;
  sushi_run_0[9][30] = 2'b01;
  sushi_run_0[9][31] = 2'b01;
  sushi_run_0[9][32] = 2'b00;
  sushi_run_0[10][0] = 2'b00;
  sushi_run_0[10][1] = 2'b00;
  sushi_run_0[10][2] = 2'b01;
  sushi_run_0[10][3] = 2'b11;
  sushi_run_0[10][4] = 2'b11;
  sushi_run_0[10][5] = 2'b10;
  sushi_run_0[10][6] = 2'b10;
  sushi_run_0[10][7] = 2'b10;
  sushi_run_0[10][8] = 2'b11;
  sushi_run_0[10][9] = 2'b10;
  sushi_run_0[10][10] = 2'b10;
  sushi_run_0[10][11] = 2'b10;
  sushi_run_0[10][12] = 2'b10;
  sushi_run_0[10][13] = 2'b10;
  sushi_run_0[10][14] = 2'b10;
  sushi_run_0[10][15] = 2'b10;
  sushi_run_0[10][16] = 2'b10;
  sushi_run_0[10][17] = 2'b10;
  sushi_run_0[10][18] = 2'b10;
  sushi_run_0[10][19] = 2'b10;
  sushi_run_0[10][20] = 2'b10;
  sushi_run_0[10][21] = 2'b10;
  sushi_run_0[10][22] = 2'b10;
  sushi_run_0[10][23] = 2'b10;
  sushi_run_0[10][24] = 2'b11;
  sushi_run_0[10][25] = 2'b10;
  sushi_run_0[10][26] = 2'b01;
  sushi_run_0[10][27] = 2'b01;
  sushi_run_0[10][28] = 2'b01;
  sushi_run_0[10][29] = 2'b01;
  sushi_run_0[10][30] = 2'b01;
  sushi_run_0[10][31] = 2'b00;
  sushi_run_0[10][32] = 2'b00;
  sushi_run_0[11][0] = 2'b00;
  sushi_run_0[11][1] = 2'b00;
  sushi_run_0[11][2] = 2'b01;
  sushi_run_0[11][3] = 2'b01;
  sushi_run_0[11][4] = 2'b11;
  sushi_run_0[11][5] = 2'b10;
  sushi_run_0[11][6] = 2'b11;
  sushi_run_0[11][7] = 2'b10;
  sushi_run_0[11][8] = 2'b10;
  sushi_run_0[11][9] = 2'b10;
  sushi_run_0[11][10] = 2'b10;
  sushi_run_0[11][11] = 2'b10;
  sushi_run_0[11][12] = 2'b10;
  sushi_run_0[11][13] = 2'b10;
  sushi_run_0[11][14] = 2'b10;
  sushi_run_0[11][15] = 2'b10;
  sushi_run_0[11][16] = 2'b10;
  sushi_run_0[11][17] = 2'b10;
  sushi_run_0[11][18] = 2'b10;
  sushi_run_0[11][19] = 2'b10;
  sushi_run_0[11][20] = 2'b11;
  sushi_run_0[11][21] = 2'b10;
  sushi_run_0[11][22] = 2'b10;
  sushi_run_0[11][23] = 2'b10;
  sushi_run_0[11][24] = 2'b10;
  sushi_run_0[11][25] = 2'b01;
  sushi_run_0[11][26] = 2'b01;
  sushi_run_0[11][27] = 2'b00;
  sushi_run_0[11][28] = 2'b00;
  sushi_run_0[11][29] = 2'b00;
  sushi_run_0[11][30] = 2'b00;
  sushi_run_0[11][31] = 2'b00;
  sushi_run_0[11][32] = 2'b00;
  sushi_run_0[12][0] = 2'b00;
  sushi_run_0[12][1] = 2'b00;
  sushi_run_0[12][2] = 2'b00;
  sushi_run_0[12][3] = 2'b01;
  sushi_run_0[12][4] = 2'b01;
  sushi_run_0[12][5] = 2'b01;
  sushi_run_0[12][6] = 2'b10;
  sushi_run_0[12][7] = 2'b10;
  sushi_run_0[12][8] = 2'b10;
  sushi_run_0[12][9] = 2'b10;
  sushi_run_0[12][10] = 2'b10;
  sushi_run_0[12][11] = 2'b10;
  sushi_run_0[12][12] = 2'b10;
  sushi_run_0[12][13] = 2'b10;
  sushi_run_0[12][14] = 2'b10;
  sushi_run_0[12][15] = 2'b10;
  sushi_run_0[12][16] = 2'b10;
  sushi_run_0[12][17] = 2'b10;
  sushi_run_0[12][18] = 2'b10;
  sushi_run_0[12][19] = 2'b10;
  sushi_run_0[12][20] = 2'b10;
  sushi_run_0[12][21] = 2'b10;
  sushi_run_0[12][22] = 2'b10;
  sushi_run_0[12][23] = 2'b10;
  sushi_run_0[12][24] = 2'b10;
  sushi_run_0[12][25] = 2'b01;
  sushi_run_0[12][26] = 2'b01;
  sushi_run_0[12][27] = 2'b00;
  sushi_run_0[12][28] = 2'b00;
  sushi_run_0[12][29] = 2'b00;
  sushi_run_0[12][30] = 2'b00;
  sushi_run_0[12][31] = 2'b00;
  sushi_run_0[12][32] = 2'b00;
  sushi_run_0[13][0] = 2'b00;
  sushi_run_0[13][1] = 2'b00;
  sushi_run_0[13][2] = 2'b00;
  sushi_run_0[13][3] = 2'b00;
  sushi_run_0[13][4] = 2'b01;
  sushi_run_0[13][5] = 2'b01;
  sushi_run_0[13][6] = 2'b10;
  sushi_run_0[13][7] = 2'b11;
  sushi_run_0[13][8] = 2'b10;
  sushi_run_0[13][9] = 2'b10;
  sushi_run_0[13][10] = 2'b10;
  sushi_run_0[13][11] = 2'b10;
  sushi_run_0[13][12] = 2'b10;
  sushi_run_0[13][13] = 2'b10;
  sushi_run_0[13][14] = 2'b10;
  sushi_run_0[13][15] = 2'b10;
  sushi_run_0[13][16] = 2'b10;
  sushi_run_0[13][17] = 2'b10;
  sushi_run_0[13][18] = 2'b10;
  sushi_run_0[13][19] = 2'b10;
  sushi_run_0[13][20] = 2'b10;
  sushi_run_0[13][21] = 2'b10;
  sushi_run_0[13][22] = 2'b10;
  sushi_run_0[13][23] = 2'b10;
  sushi_run_0[13][24] = 2'b10;
  sushi_run_0[13][25] = 2'b10;
  sushi_run_0[13][26] = 2'b01;
  sushi_run_0[13][27] = 2'b00;
  sushi_run_0[13][28] = 2'b00;
  sushi_run_0[13][29] = 2'b00;
  sushi_run_0[13][30] = 2'b00;
  sushi_run_0[13][31] = 2'b00;
  sushi_run_0[13][32] = 2'b00;
  sushi_run_0[14][0] = 2'b00;
  sushi_run_0[14][1] = 2'b00;
  sushi_run_0[14][2] = 2'b01;
  sushi_run_0[14][3] = 2'b01;
  sushi_run_0[14][4] = 2'b01;
  sushi_run_0[14][5] = 2'b11;
  sushi_run_0[14][6] = 2'b10;
  sushi_run_0[14][7] = 2'b01;
  sushi_run_0[14][8] = 2'b01;
  sushi_run_0[14][9] = 2'b11;
  sushi_run_0[14][10] = 2'b10;
  sushi_run_0[14][11] = 2'b10;
  sushi_run_0[14][12] = 2'b10;
  sushi_run_0[14][13] = 2'b10;
  sushi_run_0[14][14] = 2'b10;
  sushi_run_0[14][15] = 2'b10;
  sushi_run_0[14][16] = 2'b10;
  sushi_run_0[14][17] = 2'b10;
  sushi_run_0[14][18] = 2'b10;
  sushi_run_0[14][19] = 2'b10;
  sushi_run_0[14][20] = 2'b10;
  sushi_run_0[14][21] = 2'b10;
  sushi_run_0[14][22] = 2'b11;
  sushi_run_0[14][23] = 2'b10;
  sushi_run_0[14][24] = 2'b10;
  sushi_run_0[14][25] = 2'b10;
  sushi_run_0[14][26] = 2'b01;
  sushi_run_0[14][27] = 2'b01;
  sushi_run_0[14][28] = 2'b01;
  sushi_run_0[14][29] = 2'b00;
  sushi_run_0[14][30] = 2'b00;
  sushi_run_0[14][31] = 2'b00;
  sushi_run_0[14][32] = 2'b00;
  sushi_run_0[15][0] = 2'b00;
  sushi_run_0[15][1] = 2'b01;
  sushi_run_0[15][2] = 2'b01;
  sushi_run_0[15][3] = 2'b11;
  sushi_run_0[15][4] = 2'b10;
  sushi_run_0[15][5] = 2'b01;
  sushi_run_0[15][6] = 2'b01;
  sushi_run_0[15][7] = 2'b01;
  sushi_run_0[15][8] = 2'b01;
  sushi_run_0[15][9] = 2'b01;
  sushi_run_0[15][10] = 2'b01;
  sushi_run_0[15][11] = 2'b01;
  sushi_run_0[15][12] = 2'b10;
  sushi_run_0[15][13] = 2'b10;
  sushi_run_0[15][14] = 2'b10;
  sushi_run_0[15][15] = 2'b01;
  sushi_run_0[15][16] = 2'b10;
  sushi_run_0[15][17] = 2'b01;
  sushi_run_0[15][18] = 2'b01;
  sushi_run_0[15][19] = 2'b01;
  sushi_run_0[15][20] = 2'b10;
  sushi_run_0[15][21] = 2'b10;
  sushi_run_0[15][22] = 2'b11;
  sushi_run_0[15][23] = 2'b11;
  sushi_run_0[15][24] = 2'b10;
  sushi_run_0[15][25] = 2'b10;
  sushi_run_0[15][26] = 2'b10;
  sushi_run_0[15][27] = 2'b10;
  sushi_run_0[15][28] = 2'b01;
  sushi_run_0[15][29] = 2'b01;
  sushi_run_0[15][30] = 2'b01;
  sushi_run_0[15][31] = 2'b00;
  sushi_run_0[15][32] = 2'b00;
  sushi_run_0[16][0] = 2'b00;
  sushi_run_0[16][1] = 2'b01;
  sushi_run_0[16][2] = 2'b01;
  sushi_run_0[16][3] = 2'b01;
  sushi_run_0[16][4] = 2'b01;
  sushi_run_0[16][5] = 2'b01;
  sushi_run_0[16][6] = 2'b10;
  sushi_run_0[16][7] = 2'b10;
  sushi_run_0[16][8] = 2'b01;
  sushi_run_0[16][9] = 2'b01;
  sushi_run_0[16][10] = 2'b00;
  sushi_run_0[16][11] = 2'b01;
  sushi_run_0[16][12] = 2'b01;
  sushi_run_0[16][13] = 2'b01;
  sushi_run_0[16][14] = 2'b01;
  sushi_run_0[16][15] = 2'b01;
  sushi_run_0[16][16] = 2'b01;
  sushi_run_0[16][17] = 2'b01;
  sushi_run_0[16][18] = 2'b01;
  sushi_run_0[16][19] = 2'b01;
  sushi_run_0[16][20] = 2'b01;
  sushi_run_0[16][21] = 2'b01;
  sushi_run_0[16][22] = 2'b01;
  sushi_run_0[16][23] = 2'b01;
  sushi_run_0[16][24] = 2'b01;
  sushi_run_0[16][25] = 2'b01;
  sushi_run_0[16][26] = 2'b10;
  sushi_run_0[16][27] = 2'b10;
  sushi_run_0[16][28] = 2'b10;
  sushi_run_0[16][29] = 2'b01;
  sushi_run_0[16][30] = 2'b01;
  sushi_run_0[16][31] = 2'b00;
  sushi_run_0[16][32] = 2'b00;
  sushi_run_0[17][0] = 2'b00;
  sushi_run_0[17][1] = 2'b00;
  sushi_run_0[17][2] = 2'b00;
  sushi_run_0[17][3] = 2'b01;
  sushi_run_0[17][4] = 2'b01;
  sushi_run_0[17][5] = 2'b01;
  sushi_run_0[17][6] = 2'b01;
  sushi_run_0[17][7] = 2'b01;
  sushi_run_0[17][8] = 2'b01;
  sushi_run_0[17][9] = 2'b00;
  sushi_run_0[17][10] = 2'b00;
  sushi_run_0[17][11] = 2'b00;
  sushi_run_0[17][12] = 2'b00;
  sushi_run_0[17][13] = 2'b00;
  sushi_run_0[17][14] = 2'b00;
  sushi_run_0[17][15] = 2'b00;
  sushi_run_0[17][16] = 2'b00;
  sushi_run_0[17][17] = 2'b00;
  sushi_run_0[17][18] = 2'b00;
  sushi_run_0[17][19] = 2'b00;
  sushi_run_0[17][20] = 2'b00;
  sushi_run_0[17][21] = 2'b00;
  sushi_run_0[17][22] = 2'b00;
  sushi_run_0[17][23] = 2'b00;
  sushi_run_0[17][24] = 2'b00;
  sushi_run_0[17][25] = 2'b01;
  sushi_run_0[17][26] = 2'b01;
  sushi_run_0[17][27] = 2'b01;
  sushi_run_0[17][28] = 2'b01;
  sushi_run_0[17][29] = 2'b01;
  sushi_run_0[17][30] = 2'b00;
  sushi_run_0[17][31] = 2'b00;
  sushi_run_0[17][32] = 2'b00;
  sushi_run_0[18][0] = 2'b00;
  sushi_run_0[18][1] = 2'b00;
  sushi_run_0[18][2] = 2'b00;
  sushi_run_0[18][3] = 2'b00;
  sushi_run_0[18][4] = 2'b00;
  sushi_run_0[18][5] = 2'b00;
  sushi_run_0[18][6] = 2'b00;
  sushi_run_0[18][7] = 2'b00;
  sushi_run_0[18][8] = 2'b00;
  sushi_run_0[18][9] = 2'b00;
  sushi_run_0[18][10] = 2'b00;
  sushi_run_0[18][11] = 2'b00;
  sushi_run_0[18][12] = 2'b00;
  sushi_run_0[18][13] = 2'b00;
  sushi_run_0[18][14] = 2'b00;
  sushi_run_0[18][15] = 2'b00;
  sushi_run_0[18][16] = 2'b00;
  sushi_run_0[18][17] = 2'b00;
  sushi_run_0[18][18] = 2'b00;
  sushi_run_0[18][19] = 2'b00;
  sushi_run_0[18][20] = 2'b00;
  sushi_run_0[18][21] = 2'b00;
  sushi_run_0[18][22] = 2'b00;
  sushi_run_0[18][23] = 2'b00;
  sushi_run_0[18][24] = 2'b00;
  sushi_run_0[18][25] = 2'b00;
  sushi_run_0[18][26] = 2'b00;
  sushi_run_0[18][27] = 2'b00;
  sushi_run_0[18][28] = 2'b00;
  sushi_run_0[18][29] = 2'b00;
  sushi_run_0[18][30] = 2'b00;
  sushi_run_0[18][31] = 2'b00;
  sushi_run_0[18][32] = 2'b00;
  end

  reg [1:0] sushi_run_1 [18:0] [32:0]; //33x19 sprite [y][x]

  always @(*) begin
  sushi_run_1[0][0] = 2'b00;
  sushi_run_1[0][1] = 2'b00;
  sushi_run_1[0][2] = 2'b00;
  sushi_run_1[0][3] = 2'b00;
  sushi_run_1[0][4] = 2'b00;
  sushi_run_1[0][5] = 2'b00;
  sushi_run_1[0][6] = 2'b00;
  sushi_run_1[0][7] = 2'b00;
  sushi_run_1[0][8] = 2'b00;
  sushi_run_1[0][9] = 2'b00;
  sushi_run_1[0][10] = 2'b00;
  sushi_run_1[0][11] = 2'b00;
  sushi_run_1[0][12] = 2'b00;
  sushi_run_1[0][13] = 2'b00;
  sushi_run_1[0][14] = 2'b00;
  sushi_run_1[0][15] = 2'b00;
  sushi_run_1[0][16] = 2'b00;
  sushi_run_1[0][17] = 2'b00;
  sushi_run_1[0][18] = 2'b00;
  sushi_run_1[0][19] = 2'b00;
  sushi_run_1[0][20] = 2'b00;
  sushi_run_1[0][21] = 2'b00;
  sushi_run_1[0][22] = 2'b01;
  sushi_run_1[0][23] = 2'b01;
  sushi_run_1[0][24] = 2'b01;
  sushi_run_1[0][25] = 2'b01;
  sushi_run_1[0][26] = 2'b01;
  sushi_run_1[0][27] = 2'b01;
  sushi_run_1[0][28] = 2'b00;
  sushi_run_1[0][29] = 2'b00;
  sushi_run_1[0][30] = 2'b00;
  sushi_run_1[0][31] = 2'b00;
  sushi_run_1[0][32] = 2'b00;
  sushi_run_1[1][0] = 2'b00;
  sushi_run_1[1][1] = 2'b00;
  sushi_run_1[1][2] = 2'b00;
  sushi_run_1[1][3] = 2'b00;
  sushi_run_1[1][4] = 2'b00;
  sushi_run_1[1][5] = 2'b00;
  sushi_run_1[1][6] = 2'b00;
  sushi_run_1[1][7] = 2'b00;
  sushi_run_1[1][8] = 2'b00;
  sushi_run_1[1][9] = 2'b00;
  sushi_run_1[1][10] = 2'b00;
  sushi_run_1[1][11] = 2'b00;
  sushi_run_1[1][12] = 2'b00;
  sushi_run_1[1][13] = 2'b00;
  sushi_run_1[1][14] = 2'b00;
  sushi_run_1[1][15] = 2'b00;
  sushi_run_1[1][16] = 2'b00;
  sushi_run_1[1][17] = 2'b00;
  sushi_run_1[1][18] = 2'b00;
  sushi_run_1[1][19] = 2'b00;
  sushi_run_1[1][20] = 2'b00;
  sushi_run_1[1][21] = 2'b01;
  sushi_run_1[1][22] = 2'b01;
  sushi_run_1[1][23] = 2'b11;
  sushi_run_1[1][24] = 2'b10;
  sushi_run_1[1][25] = 2'b10;
  sushi_run_1[1][26] = 2'b10;
  sushi_run_1[1][27] = 2'b01;
  sushi_run_1[1][28] = 2'b01;
  sushi_run_1[1][29] = 2'b00;
  sushi_run_1[1][30] = 2'b00;
  sushi_run_1[1][31] = 2'b00;
  sushi_run_1[1][32] = 2'b00;
  sushi_run_1[2][0] = 2'b00;
  sushi_run_1[2][1] = 2'b00;
  sushi_run_1[2][2] = 2'b00;
  sushi_run_1[2][3] = 2'b00;
  sushi_run_1[2][4] = 2'b00;
  sushi_run_1[2][5] = 2'b00;
  sushi_run_1[2][6] = 2'b00;
  sushi_run_1[2][7] = 2'b00;
  sushi_run_1[2][8] = 2'b00;
  sushi_run_1[2][9] = 2'b00;
  sushi_run_1[2][10] = 2'b00;
  sushi_run_1[2][11] = 2'b00;
  sushi_run_1[2][12] = 2'b00;
  sushi_run_1[2][13] = 2'b00;
  sushi_run_1[2][14] = 2'b00;
  sushi_run_1[2][15] = 2'b00;
  sushi_run_1[2][16] = 2'b00;
  sushi_run_1[2][17] = 2'b00;
  sushi_run_1[2][18] = 2'b00;
  sushi_run_1[2][19] = 2'b00;
  sushi_run_1[2][20] = 2'b01;
  sushi_run_1[2][21] = 2'b01;
  sushi_run_1[2][22] = 2'b11;
  sushi_run_1[2][23] = 2'b10;
  sushi_run_1[2][24] = 2'b10;
  sushi_run_1[2][25] = 2'b10;
  sushi_run_1[2][26] = 2'b10;
  sushi_run_1[2][27] = 2'b10;
  sushi_run_1[2][28] = 2'b01;
  sushi_run_1[2][29] = 2'b01;
  sushi_run_1[2][30] = 2'b00;
  sushi_run_1[2][31] = 2'b00;
  sushi_run_1[2][32] = 2'b00;
  sushi_run_1[3][0] = 2'b00;
  sushi_run_1[3][1] = 2'b00;
  sushi_run_1[3][2] = 2'b00;
  sushi_run_1[3][3] = 2'b00;
  sushi_run_1[3][4] = 2'b00;
  sushi_run_1[3][5] = 2'b00;
  sushi_run_1[3][6] = 2'b00;
  sushi_run_1[3][7] = 2'b00;
  sushi_run_1[3][8] = 2'b00;
  sushi_run_1[3][9] = 2'b00;
  sushi_run_1[3][10] = 2'b00;
  sushi_run_1[3][11] = 2'b00;
  sushi_run_1[3][12] = 2'b00;
  sushi_run_1[3][13] = 2'b00;
  sushi_run_1[3][14] = 2'b00;
  sushi_run_1[3][15] = 2'b00;
  sushi_run_1[3][16] = 2'b00;
  sushi_run_1[3][17] = 2'b00;
  sushi_run_1[3][18] = 2'b00;
  sushi_run_1[3][19] = 2'b00;
  sushi_run_1[3][20] = 2'b01;
  sushi_run_1[3][21] = 2'b11;
  sushi_run_1[3][22] = 2'b10;
  sushi_run_1[3][23] = 2'b10;
  sushi_run_1[3][24] = 2'b10;
  sushi_run_1[3][25] = 2'b10;
  sushi_run_1[3][26] = 2'b10;
  sushi_run_1[3][27] = 2'b10;
  sushi_run_1[3][28] = 2'b10;
  sushi_run_1[3][29] = 2'b01;
  sushi_run_1[3][30] = 2'b00;
  sushi_run_1[3][31] = 2'b00;
  sushi_run_1[3][32] = 2'b00;
  sushi_run_1[4][0] = 2'b01;
  sushi_run_1[4][1] = 2'b01;
  sushi_run_1[4][2] = 2'b00;
  sushi_run_1[4][3] = 2'b00;
  sushi_run_1[4][4] = 2'b00;
  sushi_run_1[4][5] = 2'b00;
  sushi_run_1[4][6] = 2'b00;
  sushi_run_1[4][7] = 2'b00;
  sushi_run_1[4][8] = 2'b00;
  sushi_run_1[4][9] = 2'b00;
  sushi_run_1[4][10] = 2'b00;
  sushi_run_1[4][11] = 2'b00;
  sushi_run_1[4][12] = 2'b00;
  sushi_run_1[4][13] = 2'b00;
  sushi_run_1[4][14] = 2'b00;
  sushi_run_1[4][15] = 2'b00;
  sushi_run_1[4][16] = 2'b00;
  sushi_run_1[4][17] = 2'b00;
  sushi_run_1[4][18] = 2'b01;
  sushi_run_1[4][19] = 2'b01;
  sushi_run_1[4][20] = 2'b11;
  sushi_run_1[4][21] = 2'b10;
  sushi_run_1[4][22] = 2'b10;
  sushi_run_1[4][23] = 2'b10;
  sushi_run_1[4][24] = 2'b10;
  sushi_run_1[4][25] = 2'b10;
  sushi_run_1[4][26] = 2'b01;
  sushi_run_1[4][27] = 2'b01;
  sushi_run_1[4][28] = 2'b10;
  sushi_run_1[4][29] = 2'b01;
  sushi_run_1[4][30] = 2'b01;
  sushi_run_1[4][31] = 2'b00;
  sushi_run_1[4][32] = 2'b00;
  sushi_run_1[5][0] = 2'b01;
  sushi_run_1[5][1] = 2'b01;
  sushi_run_1[5][2] = 2'b01;
  sushi_run_1[5][3] = 2'b00;
  sushi_run_1[5][4] = 2'b00;
  sushi_run_1[5][5] = 2'b00;
  sushi_run_1[5][6] = 2'b00;
  sushi_run_1[5][7] = 2'b00;
  sushi_run_1[5][8] = 2'b00;
  sushi_run_1[5][9] = 2'b00;
  sushi_run_1[5][10] = 2'b00;
  sushi_run_1[5][11] = 2'b00;
  sushi_run_1[5][12] = 2'b00;
  sushi_run_1[5][13] = 2'b00;
  sushi_run_1[5][14] = 2'b00;
  sushi_run_1[5][15] = 2'b00;
  sushi_run_1[5][16] = 2'b00;
  sushi_run_1[5][17] = 2'b00;
  sushi_run_1[5][18] = 2'b01;
  sushi_run_1[5][19] = 2'b11;
  sushi_run_1[5][20] = 2'b11;
  sushi_run_1[5][21] = 2'b10;
  sushi_run_1[5][22] = 2'b10;
  sushi_run_1[5][23] = 2'b10;
  sushi_run_1[5][24] = 2'b10;
  sushi_run_1[5][25] = 2'b10;
  sushi_run_1[5][26] = 2'b10;
  sushi_run_1[5][27] = 2'b01;
  sushi_run_1[5][28] = 2'b01;
  sushi_run_1[5][29] = 2'b10;
  sushi_run_1[5][30] = 2'b01;
  sushi_run_1[5][31] = 2'b00;
  sushi_run_1[5][32] = 2'b00;
  sushi_run_1[6][0] = 2'b01;
  sushi_run_1[6][1] = 2'b01;
  sushi_run_1[6][2] = 2'b01;
  sushi_run_1[6][3] = 2'b01;
  sushi_run_1[6][4] = 2'b00;
  sushi_run_1[6][5] = 2'b00;
  sushi_run_1[6][6] = 2'b00;
  sushi_run_1[6][7] = 2'b00;
  sushi_run_1[6][8] = 2'b00;
  sushi_run_1[6][9] = 2'b00;
  sushi_run_1[6][10] = 2'b00;
  sushi_run_1[6][11] = 2'b00;
  sushi_run_1[6][12] = 2'b00;
  sushi_run_1[6][13] = 2'b00;
  sushi_run_1[6][14] = 2'b00;
  sushi_run_1[6][15] = 2'b00;
  sushi_run_1[6][16] = 2'b00;
  sushi_run_1[6][17] = 2'b00;
  sushi_run_1[6][18] = 2'b01;
  sushi_run_1[6][19] = 2'b11;
  sushi_run_1[6][20] = 2'b10;
  sushi_run_1[6][21] = 2'b10;
  sushi_run_1[6][22] = 2'b10;
  sushi_run_1[6][23] = 2'b10;
  sushi_run_1[6][24] = 2'b01;
  sushi_run_1[6][25] = 2'b10;
  sushi_run_1[6][26] = 2'b10;
  sushi_run_1[6][27] = 2'b01;
  sushi_run_1[6][28] = 2'b01;
  sushi_run_1[6][29] = 2'b10;
  sushi_run_1[6][30] = 2'b01;
  sushi_run_1[6][31] = 2'b01;
  sushi_run_1[6][32] = 2'b01;
  sushi_run_1[7][0] = 2'b00;
  sushi_run_1[7][1] = 2'b01;
  sushi_run_1[7][2] = 2'b10;
  sushi_run_1[7][3] = 2'b01;
  sushi_run_1[7][4] = 2'b00;
  sushi_run_1[7][5] = 2'b00;
  sushi_run_1[7][6] = 2'b00;
  sushi_run_1[7][7] = 2'b00;
  sushi_run_1[7][8] = 2'b00;
  sushi_run_1[7][9] = 2'b00;
  sushi_run_1[7][10] = 2'b00;
  sushi_run_1[7][11] = 2'b00;
  sushi_run_1[7][12] = 2'b00;
  sushi_run_1[7][13] = 2'b00;
  sushi_run_1[7][14] = 2'b00;
  sushi_run_1[7][15] = 2'b01;
  sushi_run_1[7][16] = 2'b01;
  sushi_run_1[7][17] = 2'b01;
  sushi_run_1[7][18] = 2'b01;
  sushi_run_1[7][19] = 2'b11;
  sushi_run_1[7][20] = 2'b10;
  sushi_run_1[7][21] = 2'b10;
  sushi_run_1[7][22] = 2'b10;
  sushi_run_1[7][23] = 2'b01;
  sushi_run_1[7][24] = 2'b01;
  sushi_run_1[7][25] = 2'b10;
  sushi_run_1[7][26] = 2'b10;
  sushi_run_1[7][27] = 2'b10;
  sushi_run_1[7][28] = 2'b10;
  sushi_run_1[7][29] = 2'b10;
  sushi_run_1[7][30] = 2'b10;
  sushi_run_1[7][31] = 2'b10;
  sushi_run_1[7][32] = 2'b01;
  sushi_run_1[8][0] = 2'b00;
  sushi_run_1[8][1] = 2'b01;
  sushi_run_1[8][2] = 2'b10;
  sushi_run_1[8][3] = 2'b01;
  sushi_run_1[8][4] = 2'b01;
  sushi_run_1[8][5] = 2'b01;
  sushi_run_1[8][6] = 2'b00;
  sushi_run_1[8][7] = 2'b01;
  sushi_run_1[8][8] = 2'b01;
  sushi_run_1[8][9] = 2'b01;
  sushi_run_1[8][10] = 2'b01;
  sushi_run_1[8][11] = 2'b01;
  sushi_run_1[8][12] = 2'b01;
  sushi_run_1[8][13] = 2'b01;
  sushi_run_1[8][14] = 2'b01;
  sushi_run_1[8][15] = 2'b01;
  sushi_run_1[8][16] = 2'b10;
  sushi_run_1[8][17] = 2'b11;
  sushi_run_1[8][18] = 2'b01;
  sushi_run_1[8][19] = 2'b01;
  sushi_run_1[8][20] = 2'b10;
  sushi_run_1[8][21] = 2'b10;
  sushi_run_1[8][22] = 2'b10;
  sushi_run_1[8][23] = 2'b01;
  sushi_run_1[8][24] = 2'b10;
  sushi_run_1[8][25] = 2'b10;
  sushi_run_1[8][26] = 2'b10;
  sushi_run_1[8][27] = 2'b10;
  sushi_run_1[8][28] = 2'b10;
  sushi_run_1[8][29] = 2'b10;
  sushi_run_1[8][30] = 2'b10;
  sushi_run_1[8][31] = 2'b01;
  sushi_run_1[8][32] = 2'b01;
  sushi_run_1[9][0] = 2'b00;
  sushi_run_1[9][1] = 2'b01;
  sushi_run_1[9][2] = 2'b01;
  sushi_run_1[9][3] = 2'b10;
  sushi_run_1[9][4] = 2'b10;
  sushi_run_1[9][5] = 2'b01;
  sushi_run_1[9][6] = 2'b01;
  sushi_run_1[9][7] = 2'b01;
  sushi_run_1[9][8] = 2'b10;
  sushi_run_1[9][9] = 2'b10;
  sushi_run_1[9][10] = 2'b10;
  sushi_run_1[9][11] = 2'b10;
  sushi_run_1[9][12] = 2'b10;
  sushi_run_1[9][13] = 2'b10;
  sushi_run_1[9][14] = 2'b10;
  sushi_run_1[9][15] = 2'b10;
  sushi_run_1[9][16] = 2'b10;
  sushi_run_1[9][17] = 2'b11;
  sushi_run_1[9][18] = 2'b10;
  sushi_run_1[9][19] = 2'b01;
  sushi_run_1[9][20] = 2'b01;
  sushi_run_1[9][21] = 2'b01;
  sushi_run_1[9][22] = 2'b01;
  sushi_run_1[9][23] = 2'b01;
  sushi_run_1[9][24] = 2'b10;
  sushi_run_1[9][25] = 2'b10;
  sushi_run_1[9][26] = 2'b10;
  sushi_run_1[9][27] = 2'b10;
  sushi_run_1[9][28] = 2'b10;
  sushi_run_1[9][29] = 2'b10;
  sushi_run_1[9][30] = 2'b01;
  sushi_run_1[9][31] = 2'b01;
  sushi_run_1[9][32] = 2'b00;
  sushi_run_1[10][0] = 2'b00;
  sushi_run_1[10][1] = 2'b00;
  sushi_run_1[10][2] = 2'b01;
  sushi_run_1[10][3] = 2'b11;
  sushi_run_1[10][4] = 2'b11;
  sushi_run_1[10][5] = 2'b10;
  sushi_run_1[10][6] = 2'b10;
  sushi_run_1[10][7] = 2'b10;
  sushi_run_1[10][8] = 2'b11;
  sushi_run_1[10][9] = 2'b10;
  sushi_run_1[10][10] = 2'b10;
  sushi_run_1[10][11] = 2'b10;
  sushi_run_1[10][12] = 2'b10;
  sushi_run_1[10][13] = 2'b10;
  sushi_run_1[10][14] = 2'b10;
  sushi_run_1[10][15] = 2'b10;
  sushi_run_1[10][16] = 2'b10;
  sushi_run_1[10][17] = 2'b10;
  sushi_run_1[10][18] = 2'b10;
  sushi_run_1[10][19] = 2'b10;
  sushi_run_1[10][20] = 2'b10;
  sushi_run_1[10][21] = 2'b10;
  sushi_run_1[10][22] = 2'b10;
  sushi_run_1[10][23] = 2'b10;
  sushi_run_1[10][24] = 2'b11;
  sushi_run_1[10][25] = 2'b10;
  sushi_run_1[10][26] = 2'b01;
  sushi_run_1[10][27] = 2'b01;
  sushi_run_1[10][28] = 2'b01;
  sushi_run_1[10][29] = 2'b01;
  sushi_run_1[10][30] = 2'b01;
  sushi_run_1[10][31] = 2'b00;
  sushi_run_1[10][32] = 2'b00;
  sushi_run_1[11][0] = 2'b00;
  sushi_run_1[11][1] = 2'b00;
  sushi_run_1[11][2] = 2'b01;
  sushi_run_1[11][3] = 2'b01;
  sushi_run_1[11][4] = 2'b11;
  sushi_run_1[11][5] = 2'b10;
  sushi_run_1[11][6] = 2'b11;
  sushi_run_1[11][7] = 2'b10;
  sushi_run_1[11][8] = 2'b10;
  sushi_run_1[11][9] = 2'b10;
  sushi_run_1[11][10] = 2'b10;
  sushi_run_1[11][11] = 2'b10;
  sushi_run_1[11][12] = 2'b10;
  sushi_run_1[11][13] = 2'b10;
  sushi_run_1[11][14] = 2'b10;
  sushi_run_1[11][15] = 2'b10;
  sushi_run_1[11][16] = 2'b10;
  sushi_run_1[11][17] = 2'b10;
  sushi_run_1[11][18] = 2'b10;
  sushi_run_1[11][19] = 2'b10;
  sushi_run_1[11][20] = 2'b11;
  sushi_run_1[11][21] = 2'b10;
  sushi_run_1[11][22] = 2'b10;
  sushi_run_1[11][23] = 2'b10;
  sushi_run_1[11][24] = 2'b10;
  sushi_run_1[11][25] = 2'b01;
  sushi_run_1[11][26] = 2'b01;
  sushi_run_1[11][27] = 2'b00;
  sushi_run_1[11][28] = 2'b00;
  sushi_run_1[11][29] = 2'b00;
  sushi_run_1[11][30] = 2'b00;
  sushi_run_1[11][31] = 2'b00;
  sushi_run_1[11][32] = 2'b00;
  sushi_run_1[12][0] = 2'b00;
  sushi_run_1[12][1] = 2'b00;
  sushi_run_1[12][2] = 2'b00;
  sushi_run_1[12][3] = 2'b01;
  sushi_run_1[12][4] = 2'b01;
  sushi_run_1[12][5] = 2'b01;
  sushi_run_1[12][6] = 2'b10;
  sushi_run_1[12][7] = 2'b10;
  sushi_run_1[12][8] = 2'b10;
  sushi_run_1[12][9] = 2'b10;
  sushi_run_1[12][10] = 2'b10;
  sushi_run_1[12][11] = 2'b10;
  sushi_run_1[12][12] = 2'b10;
  sushi_run_1[12][13] = 2'b10;
  sushi_run_1[12][14] = 2'b10;
  sushi_run_1[12][15] = 2'b10;
  sushi_run_1[12][16] = 2'b10;
  sushi_run_1[12][17] = 2'b10;
  sushi_run_1[12][18] = 2'b10;
  sushi_run_1[12][19] = 2'b10;
  sushi_run_1[12][20] = 2'b10;
  sushi_run_1[12][21] = 2'b10;
  sushi_run_1[12][22] = 2'b10;
  sushi_run_1[12][23] = 2'b10;
  sushi_run_1[12][24] = 2'b10;
  sushi_run_1[12][25] = 2'b01;
  sushi_run_1[12][26] = 2'b01;
  sushi_run_1[12][27] = 2'b00;
  sushi_run_1[12][28] = 2'b00;
  sushi_run_1[12][29] = 2'b00;
  sushi_run_1[12][30] = 2'b00;
  sushi_run_1[12][31] = 2'b00;
  sushi_run_1[12][32] = 2'b00;
  sushi_run_1[13][0] = 2'b00;
  sushi_run_1[13][1] = 2'b00;
  sushi_run_1[13][2] = 2'b00;
  sushi_run_1[13][3] = 2'b00;
  sushi_run_1[13][4] = 2'b00;
  sushi_run_1[13][5] = 2'b01;
  sushi_run_1[13][6] = 2'b01;
  sushi_run_1[13][7] = 2'b01;
  sushi_run_1[13][8] = 2'b10;
  sushi_run_1[13][9] = 2'b10;
  sushi_run_1[13][10] = 2'b10;
  sushi_run_1[13][11] = 2'b10;
  sushi_run_1[13][12] = 2'b10;
  sushi_run_1[13][13] = 2'b10;
  sushi_run_1[13][14] = 2'b10;
  sushi_run_1[13][15] = 2'b10;
  sushi_run_1[13][16] = 2'b10;
  sushi_run_1[13][17] = 2'b10;
  sushi_run_1[13][18] = 2'b10;
  sushi_run_1[13][19] = 2'b10;
  sushi_run_1[13][20] = 2'b10;
  sushi_run_1[13][21] = 2'b10;
  sushi_run_1[13][22] = 2'b10;
  sushi_run_1[13][23] = 2'b10;
  sushi_run_1[13][24] = 2'b10;
  sushi_run_1[13][25] = 2'b01;
  sushi_run_1[13][26] = 2'b00;
  sushi_run_1[13][27] = 2'b00;
  sushi_run_1[13][28] = 2'b00;
  sushi_run_1[13][29] = 2'b00;
  sushi_run_1[13][30] = 2'b00;
  sushi_run_1[13][31] = 2'b00;
  sushi_run_1[13][32] = 2'b00;
  sushi_run_1[14][0] = 2'b00;
  sushi_run_1[14][1] = 2'b00;
  sushi_run_1[14][2] = 2'b00;
  sushi_run_1[14][3] = 2'b00;
  sushi_run_1[14][4] = 2'b00;
  sushi_run_1[14][5] = 2'b00;
  sushi_run_1[14][6] = 2'b00;
  sushi_run_1[14][7] = 2'b01;
  sushi_run_1[14][8] = 2'b01;
  sushi_run_1[14][9] = 2'b01;
  sushi_run_1[14][10] = 2'b10;
  sushi_run_1[14][11] = 2'b01;
  sushi_run_1[14][12] = 2'b01;
  sushi_run_1[14][13] = 2'b11;
  sushi_run_1[14][14] = 2'b11;
  sushi_run_1[14][15] = 2'b11;
  sushi_run_1[14][16] = 2'b11;
  sushi_run_1[14][17] = 2'b10;
  sushi_run_1[14][18] = 2'b10;
  sushi_run_1[14][19] = 2'b10;
  sushi_run_1[14][20] = 2'b10;
  sushi_run_1[14][21] = 2'b10;
  sushi_run_1[14][22] = 2'b10;
  sushi_run_1[14][23] = 2'b10;
  sushi_run_1[14][24] = 2'b01;
  sushi_run_1[14][25] = 2'b01;
  sushi_run_1[14][26] = 2'b00;
  sushi_run_1[14][27] = 2'b00;
  sushi_run_1[14][28] = 2'b00;
  sushi_run_1[14][29] = 2'b00;
  sushi_run_1[14][30] = 2'b00;
  sushi_run_1[14][31] = 2'b00;
  sushi_run_1[14][32] = 2'b00;
  sushi_run_1[15][0] = 2'b00;
  sushi_run_1[15][1] = 2'b00;
  sushi_run_1[15][2] = 2'b00;
  sushi_run_1[15][3] = 2'b00;
  sushi_run_1[15][4] = 2'b00;
  sushi_run_1[15][5] = 2'b00;
  sushi_run_1[15][6] = 2'b00;
  sushi_run_1[15][7] = 2'b00;
  sushi_run_1[15][8] = 2'b01;
  sushi_run_1[15][9] = 2'b11;
  sushi_run_1[15][10] = 2'b10;
  sushi_run_1[15][11] = 2'b10;
  sushi_run_1[15][12] = 2'b01;
  sushi_run_1[15][13] = 2'b01;
  sushi_run_1[15][14] = 2'b01;
  sushi_run_1[15][15] = 2'b01;
  sushi_run_1[15][16] = 2'b01;
  sushi_run_1[15][17] = 2'b11;
  sushi_run_1[15][18] = 2'b10;
  sushi_run_1[15][19] = 2'b10;
  sushi_run_1[15][20] = 2'b10;
  sushi_run_1[15][21] = 2'b10;
  sushi_run_1[15][22] = 2'b10;
  sushi_run_1[15][23] = 2'b10;
  sushi_run_1[15][24] = 2'b01;
  sushi_run_1[15][25] = 2'b00;
  sushi_run_1[15][26] = 2'b00;
  sushi_run_1[15][27] = 2'b00;
  sushi_run_1[15][28] = 2'b00;
  sushi_run_1[15][29] = 2'b00;
  sushi_run_1[15][30] = 2'b00;
  sushi_run_1[15][31] = 2'b00;
  sushi_run_1[15][32] = 2'b00;
  sushi_run_1[16][0] = 2'b00;
  sushi_run_1[16][1] = 2'b00;
  sushi_run_1[16][2] = 2'b00;
  sushi_run_1[16][3] = 2'b00;
  sushi_run_1[16][4] = 2'b00;
  sushi_run_1[16][5] = 2'b00;
  sushi_run_1[16][6] = 2'b00;
  sushi_run_1[16][7] = 2'b00;
  sushi_run_1[16][8] = 2'b01;
  sushi_run_1[16][9] = 2'b01;
  sushi_run_1[16][10] = 2'b01;
  sushi_run_1[16][11] = 2'b10;
  sushi_run_1[16][12] = 2'b01;
  sushi_run_1[16][13] = 2'b00;
  sushi_run_1[16][14] = 2'b00;
  sushi_run_1[16][15] = 2'b00;
  sushi_run_1[16][16] = 2'b01;
  sushi_run_1[16][17] = 2'b01;
  sushi_run_1[16][18] = 2'b01;
  sushi_run_1[16][19] = 2'b01;
  sushi_run_1[16][20] = 2'b01;
  sushi_run_1[16][21] = 2'b10;
  sushi_run_1[16][22] = 2'b10;
  sushi_run_1[16][23] = 2'b01;
  sushi_run_1[16][24] = 2'b01;
  sushi_run_1[16][25] = 2'b00;
  sushi_run_1[16][26] = 2'b00;
  sushi_run_1[16][27] = 2'b00;
  sushi_run_1[16][28] = 2'b00;
  sushi_run_1[16][29] = 2'b00;
  sushi_run_1[16][30] = 2'b00;
  sushi_run_1[16][31] = 2'b00;
  sushi_run_1[16][32] = 2'b00;
  sushi_run_1[17][0] = 2'b00;
  sushi_run_1[17][1] = 2'b00;
  sushi_run_1[17][2] = 2'b00;
  sushi_run_1[17][3] = 2'b00;
  sushi_run_1[17][4] = 2'b00;
  sushi_run_1[17][5] = 2'b00;
  sushi_run_1[17][6] = 2'b00;
  sushi_run_1[17][7] = 2'b00;
  sushi_run_1[17][8] = 2'b00;
  sushi_run_1[17][9] = 2'b00;
  sushi_run_1[17][10] = 2'b01;
  sushi_run_1[17][11] = 2'b01;
  sushi_run_1[17][12] = 2'b01;
  sushi_run_1[17][13] = 2'b00;
  sushi_run_1[17][14] = 2'b00;
  sushi_run_1[17][15] = 2'b00;
  sushi_run_1[17][16] = 2'b00;
  sushi_run_1[17][17] = 2'b00;
  sushi_run_1[17][18] = 2'b00;
  sushi_run_1[17][19] = 2'b01;
  sushi_run_1[17][20] = 2'b11;
  sushi_run_1[17][21] = 2'b10;
  sushi_run_1[17][22] = 2'b01;
  sushi_run_1[17][23] = 2'b01;
  sushi_run_1[17][24] = 2'b00;
  sushi_run_1[17][25] = 2'b00;
  sushi_run_1[17][26] = 2'b00;
  sushi_run_1[17][27] = 2'b00;
  sushi_run_1[17][28] = 2'b00;
  sushi_run_1[17][29] = 2'b00;
  sushi_run_1[17][30] = 2'b00;
  sushi_run_1[17][31] = 2'b00;
  sushi_run_1[17][32] = 2'b00;
  sushi_run_1[18][0] = 2'b00;
  sushi_run_1[18][1] = 2'b00;
  sushi_run_1[18][2] = 2'b00;
  sushi_run_1[18][3] = 2'b00;
  sushi_run_1[18][4] = 2'b00;
  sushi_run_1[18][5] = 2'b00;
  sushi_run_1[18][6] = 2'b00;
  sushi_run_1[18][7] = 2'b00;
  sushi_run_1[18][8] = 2'b00;
  sushi_run_1[18][9] = 2'b00;
  sushi_run_1[18][10] = 2'b00;
  sushi_run_1[18][11] = 2'b00;
  sushi_run_1[18][12] = 2'b00;
  sushi_run_1[18][13] = 2'b00;
  sushi_run_1[18][14] = 2'b00;
  sushi_run_1[18][15] = 2'b00;
  sushi_run_1[18][16] = 2'b00;
  sushi_run_1[18][17] = 2'b00;
  sushi_run_1[18][18] = 2'b00;
  sushi_run_1[18][19] = 2'b01;
  sushi_run_1[18][20] = 2'b01;
  sushi_run_1[18][21] = 2'b01;
  sushi_run_1[18][22] = 2'b01;
  sushi_run_1[18][23] = 2'b00;
  sushi_run_1[18][24] = 2'b00;
  sushi_run_1[18][25] = 2'b00;
  sushi_run_1[18][26] = 2'b00;
  sushi_run_1[18][27] = 2'b00;
  sushi_run_1[18][28] = 2'b00;
  sushi_run_1[18][29] = 2'b00;
  sushi_run_1[18][30] = 2'b00;
  sushi_run_1[18][31] = 2'b00;
  sushi_run_1[18][32] = 2'b00;
  end




  //unused outputs
  assign uio_out = 0;
  assign uio_oe  = 0; 



  //vga signals
  reg h_sync;
  reg v_sync;
  reg [1:0] r;
  reg [1:0] g;
  reg [1:0] b;

  reg display_on;
  reg [9:0] pix_x;
  reg [9:0] pix_y;


  //output
  assign uo_out = {h_sync, b[0], g[0], r[0], v_sync, b[1], g[1], r[1]};


  
  //hvsync gen
  always @(posedge clk) begin

        if (!rst_n) begin
            pix_x        <= 0;
            pix_y        <= 0;
            h_sync       <= 1;
            v_sync       <= 1;
        end
        else begin
            pix_x        <= (pix_x >= H_MAX) ? 0: pix_x + 1;
            pix_y        <= (pix_y >= V_MAX) ? 0: ((pix_x >= H_MAX) ? pix_y + 1 : pix_y);
            h_sync       <= (pix_x >= H_SYNC_START) && (pix_x <= H_SYNC_END);
            v_sync       <= (pix_y >= V_SYNC_START) && (pix_y <= V_SYNC_END);
        end
    end

    assign display_on = (pix_x < H_DISPLAY) && (pix_y < V_DISPLAY);



  //counter
  reg [4:0] counter;

  always @(posedge v_sync) begin
    if(!rst_n) begin
      counter <= 0;
    end
    else begin
      counter <= counter + 1;
    end
  end

  reg [9:0]sprite_x;
  reg [9:0]sprite_y;

  always @(posedge v_sync) begin
    if(!rst_n) begin
      sprite_x <= SPRITE_X_START;
      sprite_y <= SPRITE_Y_START;
    end
    else begin
      sprite_x <= sprite_x + 1;
    end
  end



  //pixel output
  reg [5:0] layer1_rgb;
  reg [5:0] sushi_0_rgb;
  reg [5:0] sushi_1_rgb;
  wire [5:0] background_rgb;

  always @(*) begin
    case(sushi_run_0[(pix_y - sprite_y) >> 3][(pix_x - sprite_x) >> 3]) 
      0: sushi_0_rgb = 6'b001100;
      1: sushi_0_rgb = 6'b000000;
      2: sushi_0_rgb = 6'b111111;
      3: sushi_0_rgb = 6'b101010;
      default: sushi_0_rgb = 6'b001100;
    endcase

    case(sushi_run_1[(pix_y - sprite_y) >> 3][(pix_x - sprite_x) >> 3]) 
      0: sushi_1_rgb = 6'b001100;
      1: sushi_1_rgb = 6'b000000;
      2: sushi_1_rgb = 6'b111111;
      3: sushi_1_rgb = 6'b101010;
      default: sushi_0_rgb = 6'b001100;
    endcase

  end

  // assign sushi_0_rgb = sushi_run_0[(pix_y - sprite_y) >> 3][(pix_x - sprite_x) >> 3];
  // assign sushi_1_rgb = sushi_run_1[(pix_y - sprite_y) >> 3][(pix_x - sprite_x) >> 3];
  assign background_rgb = {2'b01, 2'b01, 2'b10};


  always @(posedge clk) begin
    if(!rst_n) begin
      layer1_rgb <= background_rgb;
    end
    else if(//inside sprite
            display_on &&
            pix_x >= sprite_x && 
            pix_x < sprite_x + SPRITE_WIDTH &&
            pix_y >= sprite_y && 
            pix_y < sprite_y + SPRITE_HEIGHT) begin
                //bitmask
              if(counter[4]) begin
                layer1_rgb <= sushi_0_rgb == 6'b001100 ? background_rgb : sushi_0_rgb;
              end
              else begin
                layer1_rgb <= sushi_1_rgb == 6'b001100 ? background_rgb : sushi_1_rgb;
              end
    end
    else begin 
        //background color
        layer1_rgb <= background_rgb;
    end
    
  end

  always @(*)begin
      {r,g,b} = layer1_rgb;
  end

endmodule




